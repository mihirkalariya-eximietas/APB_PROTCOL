/////////////////////////////////////////////////////////////////
//  file name   : apb_define.sv
//  module name : apb DEFINE CLASS
//////////////////////////////////////////////////////////////////

`ifndef APB_DEFINES_SV
`define APB_DEFINES_SV

`define DATA_WIDTH 32 
`define ADDR_WIDTH 32
`define DEPTH 255

`endif




